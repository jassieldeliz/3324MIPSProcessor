//Written by Jassiel Deliz

`timescale 1ns/10ps
module cpu5_testbench();

reg  [31:0] instrbus;
reg  [31:0] instrbusin[0:63];
wire [31:0] iaddrbus, daddrbus;
reg  [31:0] iaddrbusout[0:63], daddrbusout[0:63];
wire [31:0] databus;
reg  [31:0] databusk, databusin[0:63], databusout[0:63];
reg         clk, reset;
reg         clkd;

reg [31:0] dontcare;
integer error, k, ntests;

	parameter Rformat	= 6'b000000;
	parameter ADDI		= 6'b000011;
	parameter SUBI		= 6'b000010;
	parameter XORI		= 6'b000001;
	parameter ANDI		= 6'b001111;
	parameter ORI		= 6'b001100;
	parameter LW		= 6'b011110;
	parameter SW		= 6'b011111;
	parameter BEQ		= 6'b110000;
	parameter BNE		= 6'b110001;
	parameter ADD		= 6'b000011;
	parameter SUB		= 6'b000010;
	parameter XOR		= 6'b000001;
	parameter AND		= 6'b000111;
	parameter OR		= 6'b000100;
	parameter SLT		= 6'b110110;
	parameter SLE		= 6'b110111;

cpu5 dut(.reset(reset),.clk(clk),.iaddrbus(iaddrbus),.ibus(instrbus),.daddrbus(daddrbus),.databus(databus));

initial begin
dontcare = 32'hx;

//* ADDI  R20, R0, #-1
iaddrbusout[0] = 32'h00000000;
//            opcode source1   dest      Immediate...
instrbusin[0]={ADDI, 5'b00000, 5'b10100, 16'h0000};

daddrbusout[0] = dontcare;
databusin[0] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[0] = dontcare;

//* ADDI  R21, R0, #1
iaddrbusout[1] = 32'h00000004;
//            opcode source1   dest      Immediate...
instrbusin[1]={ADDI, 5'b00000, 5'b10101, 16'hFFFF};

daddrbusout[1] = dontcare;
databusin[1] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[1] = dontcare;

//* SUBI  R22, R0, #2
iaddrbusout[2] = 32'h00000008;
//            opcode source1   dest      Immediate...
instrbusin[2]={SUBI, 5'b00000, 5'b10110, 16'hFF45};

daddrbusout[2] = dontcare;
databusin[2] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[2] = dontcare;

//* LW     R24, 0(R20)
iaddrbusout[3] = 32'h0000000C;
//            opcode source1   dest      Immediate...
instrbusin[3]={LW, 5'b10100, 5'b11000, 16'h00FF};

daddrbusout[3] = 32'h000000FF;
databusin[3] = 32'hCCCCCCCC;
databusout[3] = dontcare;

//* LW     R25, 0(R21)
iaddrbusout[4] = 32'h00000010;
//            opcode source1   dest      Immediate...
instrbusin[4]={LW, 5'b10101, 5'b11001, 16'hFF00};

daddrbusout[4] = 32'hFFFFFEFF;
databusin[4] = 32'hAAAAAAAA;
databusout[4] = dontcare;

//* SW     1000(R22), R20
iaddrbusout[5] = 32'h00000014;
//            opcode source1   dest      Immediate...
instrbusin[5]={SW, 5'b10110, 5'b10100, 16'h0000};

daddrbusout[5] = 32'h000000BB;
databusin[5] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[5] = 32'h00000000;

//* SW     2(R0), R21
iaddrbusout[6] = 32'h00000018;
//            opcode source1   dest      Immediate...
instrbusin[6]={SW, 5'b00000, 5'b10101, 16'h00FF};

daddrbusout[6] = 32'h000000FF;
databusin[6] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[6] = 32'hFFFFFFFF;

//* SUB   R26, R24, R25
iaddrbusout[7] = 32'h0000001C;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[7]={Rformat, 5'b11000, 5'b11001, 5'b11010, 5'b00000, SUB};

daddrbusout[7] = dontcare;
databusin[7] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[7] = dontcare;

//* XORI  R17, R24, 5564
iaddrbusout[8] = 32'h00000020;
//            opcode source1   dest      Immediate...
instrbusin[8]={XORI, 5'b11000, 5'b10001, 16'h5564};

daddrbusout[8] = dontcare;
databusin[8] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[8] = dontcare;

//* OR   R27, R24, R25
iaddrbusout[9] = 32'h00000024;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[9]={Rformat, 5'b11000, 5'b11001, 5'b11011, 5'b00000, OR};

daddrbusout[9] = dontcare;
databusin[9] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[9] = dontcare;

//* SUBI   R18, R24, F0F0             
iaddrbusout[10] = 32'h00000028;
//            opcode source1   dest      Immediate...
instrbusin[10]={SUBI, 5'b11000, 5'b10010, 16'hF0F0};

daddrbusout[10] = dontcare;
databusin[10] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[10] = dontcare;

//* XOR    R28, R24, R0           
iaddrbusout[11] = 32'h0000002C;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[11]={Rformat, 5'b11000, 5'b00000, 5'b11100, 5'b00000, XOR};

daddrbusout[11] = dontcare;
databusin[11] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[11] = dontcare;

//* ADDI   R19, R24, 3324
iaddrbusout[12] = 32'h00000030;
//            opcode source1   dest      Immediate...
instrbusin[12]={ADDI, 5'b11000, 5'b10011, 16'h3324};

daddrbusout[12] = dontcare;
databusin[12] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[12] = dontcare;

//* SUB    R29, R24, R25
iaddrbusout[13] = 32'h00000034;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[13]={Rformat, 5'b11000, 5'b11001, 5'b11101, 5'b00000, SUB};

daddrbusout[13] = dontcare;
databusin[13] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[13] = dontcare;

//* ANDI    R20, R24, 4567
iaddrbusout[14] = 32'h00000038;
//            opcode source1   dest      Immediate...
instrbusin[14]={ANDI, 5'b11000, 5'b10100, 16'h4567};

daddrbusout[14] = dontcare;
databusin[14] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[14] = dontcare;

//* ADD     R30, R24, R25
iaddrbusout[15] = 32'h0000003C;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[15]={Rformat, 5'b11000, 5'b11001, 5'b11110, 5'b00000, ADD};

daddrbusout[15] = dontcare;
databusin[15] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[15] =  dontcare;

//* SW     0(R26),  R26
iaddrbusout[16] = 32'h0000040;
//            opcode source1   dest      Immediate...
instrbusin[16]={SW, 5'b11010, 5'b11010, 16'h5574};

daddrbusout[16] = 32'h22227796;
databusin[16] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[16] = 32'h22222222;

//18* SW     0(R17),  R27
iaddrbusout[17] = 32'h0000044;
//            opcode source1   dest      Immediate...
instrbusin[17]={SW, 5'b10001, 5'b11011, 16'h0000};

daddrbusout[17] = 32'hCCCC99A8;
databusin[17] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[17] = 32'hEEEEEEEE;

//19* SW     1000(R18),  R28           
iaddrbusout[18] = 32'h00000048;
//            opcode source1   dest      Immediate...
instrbusin[18]={SW, 5'b10010, 5'b11100, 16'hFF00};

daddrbusout[18] = 32'hCCCCDADC;
databusin[18] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[18] = 32'hxxxxxxxx;

//20* SW     0(R19),  R29
iaddrbusout[19] = 32'h0000004C;
//            opcode source1   dest      Immediate...
instrbusin[19]={SW, 5'b10011, 5'b11101, 16'hAC65};

daddrbusout[19] = 32'hCCCCAC55;
databusin[19] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[19] = 32'h22222222;

//21* SW     0(R20),  R30
iaddrbusout[20] = 32'h00000050;
//            opcode source1   dest      Immediate...
instrbusin[20]={SW, 5'b10100, 5'b11110, 16'h8956};

daddrbusout[20] = 32'hFFFFCD9A;
databusin[20] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[20] = 32'h77777776;


//22* SLE  R1,  R0,  R21
iaddrbusout[21] = 32'h00000054;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[21]={Rformat, 5'b00000, 5'b10101, 5'b00001, 5'b00000, SLE};
daddrbusout[21] = dontcare;
databusin[21]   = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[21]  = dontcare;

//* XORI R5,  R0, #1
iaddrbusout[22] = 32'h00000058;
//            opcode source1   dest      Immediate...
instrbusin[22]={XORI, 5'b00000, 5'b00101, 16'h0001};
daddrbusout[22] = dontcare;
databusin[22] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[22] = dontcare;

//* SUBI R6,  R0, 0378
iaddrbusout[23] = 32'h0000005C;
//            opcode source1   dest      Immediate...
instrbusin[23]={SUBI, 5'b00000, 5'b00110, 16'h0378};
daddrbusout[23] = dontcare;
databusin[23] =   32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[23] =  dontcare;

//* BNE  R0,  R1, A001
iaddrbusout[24] = 32'h00000060;
//            opcode source1   dest      Immediate...
instrbusin[24]={BNE, 5'b00001, 5'b00000, 16'hA001};
daddrbusout[24] = dontcare;
databusin[24] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[24] = dontcare;

//* ORI R8,  R0, 5593
iaddrbusout[25] = 32'h00000064;
//            opcode source1   dest      Immediate...
instrbusin[25]={ORI, 5'b00000, 5'b01000, 16'h5593};
daddrbusout[25] = dontcare;
databusin[25] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[25] = dontcare;

//* SLE  R2,  R0, R0
iaddrbusout[26] = 32'hFFFE8068;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[26]={Rformat, 5'b00000, 5'b00000, 5'b00010, 5'b00000, SLE};
daddrbusout[26] = dontcare;
databusin[26] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[26] = dontcare;

//* NOP
iaddrbusout[27] = 32'hFFFE806C;
//                   oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[27] = 32'b00000000000000000000000000000000;
daddrbusout[27] = dontcare;
databusin[27] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[27] = dontcare;

//* NOP
iaddrbusout[28] = 32'hFFFE8070;
//                   oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[28] = 32'b00000000000000000000000000000011;
daddrbusout[28] = dontcare;
databusin[28]  = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[28] = dontcare;

//* BNE  R0,  R2, 0787
iaddrbusout[29] = 32'hFFFE8074;
//            opcode source1   dest      Immediate...
instrbusin[29]={BNE, 5'b00010, 5'b00000, 16'h0787};
daddrbusout[29] = dontcare;
databusin[29] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[29] = dontcare;

//* NOP
iaddrbusout[30] = 32'hFFFE8078;
//                   oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[30] = 32'b00000000000000000000000000000111;
daddrbusout[30] = dontcare;
databusin[30] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[30] = dontcare;

//* BEQ  R2,  R2, 5BAC
iaddrbusout[31] = 32'hFFFE9E94;
//            opcode source1   dest      Immediate...
instrbusin[31]={BEQ, 5'b00010, 5'b00010, 16'h5BAc};
daddrbusout[31] = dontcare;
databusin[31] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[31] = dontcare;

//* XORI R20, R0, 3333
iaddrbusout[32] = 32'hFFFE9E98;
//            opcode source1   dest      Immediate...
instrbusin[32]={XORI, 5'b00000, 5'b10100, 16'h3333};
daddrbusout[32] = dontcare;
databusin[32] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[32] = dontcare;

//* NOP
iaddrbusout[33] = 32'h00000D48;
//                   oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[33] = 32'b11000000000000000000000000000000;
daddrbusout[33] = dontcare;
databusin[33] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[33] = dontcare;

//* NOP
iaddrbusout[34] = 32'h00000D4C;
//                   oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[34] = 32'b00000011000000000000000000000000;
daddrbusout[34] = dontcare;
databusin[34] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[34] = dontcare;

//* NOP
iaddrbusout[35] = 32'h00000D4C;
//                   oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[35] = 32'b00000000110000000000000000000000;
daddrbusout[35] = dontcare;
databusin[35] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[35] = dontcare;

//* SUBI  R20, R0, 5546
iaddrbusout[36] = 32'h00000D50;
//            opcode source1   dest      Immediate...
instrbusin[36]={SUBI, 5'b00000, 5'b10100, 16'h5546};

daddrbusout[36] = dontcare;
databusin[36] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[36] = dontcare;

//* ADDI  R21, R0, #1
iaddrbusout[37] = 32'h00000D54;
//            opcode source1   dest      Immediate...
instrbusin[37]={ADDI, 5'b00000, 5'b10101, 16'hFFFF};

daddrbusout[37] = dontcare;
databusin[37] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[37] = dontcare;

//* ADDI  R22, R0, #2
iaddrbusout[38] = 32'h00000D58;
//            opcode source1   dest      Immediate...
instrbusin[38]={ADDI, 5'b00000, 5'b10110, 16'h0088};

daddrbusout[38] = dontcare;
databusin[38] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[38] = dontcare;

//* LW     R24, 0(R20)
iaddrbusout[39] = 32'h00000D5C;
//            opcode source1   dest      Immediate...
instrbusin[39]={LW, 5'b10100, 5'b11000, 16'h00FF};

daddrbusout[39] = 32'hFFFFABB9;
databusin[39] = 32'hCCCCCCCC;
databusout[39] = dontcare;

//* LW     R25, 0(R21)
iaddrbusout[40] = 32'h00000D60;
//            opcode source1   dest      Immediate...
instrbusin[40]={LW, 5'b10101, 5'b11001, 16'hFF00};

daddrbusout[40] = 32'hFFFFFEFF;
databusin[40] = 32'hAAAAAAAA;
databusout[40] = dontcare;

//* SW     1000(R22), R20
iaddrbusout[41] = 32'h00000D64;
//            opcode source1   dest      Immediate...
instrbusin[41]={SW, 5'b10110, 5'b10100, 16'h0000};

daddrbusout[41] = 32'h00000088;
databusin[41] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[41] = 32'hFFFFAABA;

//* SW     2(R0), R21
iaddrbusout[42] = 32'h00000D68;
//            opcode source1   dest      Immediate...
instrbusin[42]={SW, 5'b00000, 5'b10101, 16'h00FF};

daddrbusout[42] = 32'h000000FF;
databusin[42] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[42] = 32'hFFFFFFFF;

//* XOR   R26, R24, R25
iaddrbusout[43] = 32'h00000D6C;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[43]={Rformat, 5'b11000, 5'b11001, 5'b11010, 5'b00000, XOR};

daddrbusout[43] = dontcare;
databusin[43] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[43] = dontcare;

//* ANDI  R17, R24, 6420
iaddrbusout[44] = 32'h00000D70;
//            opcode source1   dest      Immediate...
instrbusin[44]={ANDI, 5'b11000, 5'b10001, 16'h6420};

daddrbusout[44] = dontcare;
databusin[44] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[44] = dontcare;

//* OR   R27, R24, R25
iaddrbusout[45] = 32'h00000D74;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[45]={Rformat, 5'b11000, 5'b11001, 5'b11011, 5'b00000, OR};

daddrbusout[45] = dontcare;
databusin[45] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[45] = dontcare;

//* SUBI   R18, R24, 5546             
iaddrbusout[46] = 32'h00000D78;
//            opcode source1   dest      Immediate...
instrbusin[46]={SUBI, 5'b11000, 5'b10010, 16'h5546};

daddrbusout[46] = dontcare;
databusin[46] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[46] = dontcare;

//* ADD    R28, R24, R0           
iaddrbusout[47] = 32'h00000D7C;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[47]={Rformat, 5'b11000, 5'b00000, 5'b11100, 5'b00000, ADD};

daddrbusout[47] = dontcare;
databusin[47] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[47] = dontcare;

//* ANDI   R19, R24, 6647
iaddrbusout[48] = 32'h00000D80;
//            opcode source1   dest      Immediate...
instrbusin[48]={ANDI, 5'b11000, 5'b10011, 16'h6647};

daddrbusout[48] = dontcare;
databusin[48] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[48] = dontcare;

//* OR    R29, R24, R25
iaddrbusout[49] = 32'h00000D84;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[49]={Rformat, 5'b11000, 5'b11001, 5'b11101, 5'b00000, OR};

daddrbusout[49] = dontcare;
databusin[49] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[49] = dontcare;

//* ADDI    R20, R24, 5680
iaddrbusout[50] = 32'h00000D88;
//            opcode source1   dest      Immediate...
instrbusin[50]={ADDI, 5'b11000, 5'b10100, 16'h5680};

daddrbusout[50] = dontcare;
databusin[50] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[50] = dontcare;

//* AND     R30, R24, R25
iaddrbusout[51] = 32'h00000D8C;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[51]={Rformat, 5'b11000, 5'b11001, 5'b11110, 5'b00000, AND};

daddrbusout[51] = dontcare;
databusin[51] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[51] =  dontcare;

//* SW     0(R26),  R26
iaddrbusout[52] = 32'h00000D90;
//            opcode source1   dest      Immediate...
instrbusin[52]={SW, 5'b11010, 5'b11010, 16'h0FF0};

daddrbusout[52] = 32'h66667656;
databusin[52] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[52] = 32'h66666666;

//* SW     0(R17),  R27
iaddrbusout[53] = 32'h00000D94;
//            opcode source1   dest      Immediate...
instrbusin[53]={SW, 5'b10001, 5'b11011, 16'hFFFF};

daddrbusout[53] = 32'h000043FF;
databusin[53] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[53] = 32'hEEEEEEEE;

//* SW     1000(R18),  R28           
iaddrbusout[54] = 32'h00000D98;
//            opcode source1   dest      Immediate...
instrbusin[54]={SW, 5'b10010, 5'b11100, 16'h8745};

daddrbusout[54] = 32'hCCCBFECB;
databusin[54] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[54] = 32'hxxxxxxxx;

//* SW     0(R19),  R29
iaddrbusout[55] = 32'h00000D9C;
//            opcode source1   dest      Immediate...
instrbusin[55]={SW, 5'b10011, 5'b11101, 16'h1123};

daddrbusout[55] = 32'h00005567;
databusin[55] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[55] = 32'hEEEEEEEE;

//* SW     0(R20),  R30
iaddrbusout[56] = 32'h00000DA0;
//            opcode source1   dest      Immediate...
instrbusin[56]={SW, 5'b10100, 5'b11110, 16'h0952};

daddrbusout[56] = 32'hCCCD2C9E;
databusin[56] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[56] = 32'h88888888;


//* SLT  R1,  R0,  R21
iaddrbusout[57] = 32'h00000DA4;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[57]={Rformat, 5'b00000, 5'b10101, 5'b00001, 5'b00000, SLT};
daddrbusout[57] = dontcare;
databusin[57]   = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[57]  = dontcare;

//* SUBI R5,  R0, #1
iaddrbusout[58] = 32'h00000DA8;
//            opcode source1   dest      Immediate...
instrbusin[58]={SUBI, 5'b00000, 5'b00101, 16'h0001};
daddrbusout[58] = dontcare;
databusin[58] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[58] = dontcare;

//* XORI R6,  R0, #1
iaddrbusout[59] = 32'h00000DAC;
//            opcode source1   dest      Immediate...
instrbusin[59]={XORI, 5'b00000, 5'b00110, 16'h0001};
daddrbusout[59] = dontcare;
databusin[59] =   32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[59] =  dontcare;

//* BEQ  R0,  R1, #10
iaddrbusout[60] = 32'h00000DB0;
//            opcode source1   dest      Immediate...
instrbusin[60]={BEQ, 5'b00001, 5'b00000, 16'h000A};
daddrbusout[60] = dontcare;
databusin[60] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[60] = dontcare;

//* ANDI R8,  R0, #1
iaddrbusout[61] = 32'h00000DB4;
//            opcode source1   dest      Immediate...
instrbusin[61]={ANDI, 5'b00000, 5'b01000, 16'h0001};
daddrbusout[61] = dontcare;
databusin[61] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[61] = dontcare;

//* SLT  R2,  R0, R0
iaddrbusout[62] = 32'h00000DB8;
//             opcode   source1   source2   dest      shift     Function...
instrbusin[62]={Rformat, 5'b00000, 5'b00000, 5'b00010, 5'b00000, SLT};
daddrbusout[62] = dontcare;
databusin[62] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[62] = dontcare;

//* NOP
iaddrbusout[63] = 32'h00000DBC;
//                   oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[63] = 32'b00000000000000000000000000000000;
daddrbusout[63] = dontcare;
databusin[63] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[63] = dontcare;

// (no. instructions) + (no. loads) + 2*(no. stores) = 70 + 4 + 2*15 = 102
ntests = 102;

$timeformat(-9,1,"ns",12);

end


//assumes positive edge FF.
//testbench reads databus when clk high, writes databus when clk low.
assign databus = clkd ? 32'bz : databusk;

//Change inputs in middle of period (falling edge).
initial begin
  error = 0;
  clkd =1;
  clk=1;
  $display ("Time=%t\n  clk=%b", $realtime, clk);
  databusk = 32'bz;

  //extended reset to set up PC MUX
  reset = 1;
  $display ("reset=%b", reset);
  #5
  clk=0;
  clkd=0;
  $display ("Time=%t\n  clk=%b", $realtime, clk);
  #5

  clk=1;
  clkd=1;
  $display ("Time=%t\n  clk=%b", $realtime, clk);
  #5
  clk=0;
  clkd=0;
  $display ("Time=%t\n  clk=%b", $realtime, clk);
  #5
  $display ("Time=%t\n  clk=%b", $realtime, clk);

for (k=0; k<= 63; k=k+1) begin
    clk=1;
    $display ("Time=%t\n  clk=%b", $realtime, clk);
    #2
    clkd=1;
    #3
    $display ("Time=%t\n  clk=%b", $realtime, clk);
    reset = 0;
    $display ("reset=%b", reset);


    //set load data for 3rd previous instruction
    if (k >=3)
      databusk = databusin[k-3];

    //check PC for this instruction
    if (k >= 0) begin
      $display ("  Testing PC for instruction %d", k);
      $display ("    Your iaddrbus =    %b", iaddrbus);
      $display ("    Correct iaddrbus = %b", iaddrbusout[k]);
      if (iaddrbusout[k] !== iaddrbus) begin
        $display ("    -------------ERROR. A Mismatch Has Occured-----------");
        error = error + 1;
      end
    end

    //put next instruction on ibus
    instrbus=instrbusin[k];
    $display ("  instrbus=%b %b %b %b %b for instruction %d:", instrbus[31:26], instrbus[25:21], instrbus[20:16], instrbus[15:11], instrbus[10:0], k);

    //check data address from 3rd previous instruction
    if ( (k >= 3) && (daddrbusout[k-3] !== dontcare) ) begin
      $display ("  Testing data address for instruction %d:", k-3);
      $display ("    Your daddrbus =    %b", daddrbus);
      $display ("    Correct daddrbus = %b", daddrbusout[k-3]);
      if (daddrbusout[k-3] !== daddrbus) begin
        $display ("    -------------ERROR. A Mismatch Has Occured-----------");
        error = error + 1;
      end
    end

    //check store data from 3rd previous instruction
    if ( (k >= 3) && (databusout[k-3] !== dontcare) ) begin
      $display ("  Testing store data for instruction %d:", k-3);
      $display ("    Your databus =    %b", databus);
      $display ("    Correct databus = %b", databusout[k-3]);
      if (databusout[k-3] !== databus) begin
        $display ("    -------------ERROR. A Mismatch Has Occured-----------");
        error = error + 1;
      end
    end

    clk = 0;
    $display ("Time=%t\n  clk=%b", $realtime, clk);
    #2
    clkd = 0;
    #3
    $display ("Time=%t\n  clk=%b", $realtime, clk);
  end

  if ( error !== 0) begin
    $display("--------- SIMULATION UNSUCCESFUL - MISMATCHES HAVE OCCURED ----------");
    $display(" No. Of Errors = %d", error);
  end
  if ( error == 0)
    $display("---------YOU DID IT!! SIMULATION SUCCESFULLY FINISHED----------");
end

endmodule
